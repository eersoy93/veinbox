/* DESCRIPTION: VeinBox simulation data types source file
 * AUTHOR: Erdem Ersoy (eersoy93)
 * See README.md for copyright and license.
 */

module simulation

type DataTypeBool                = int
type DataTypeByte                = u8
type DataTypeCChar               = i8
type DataTypeDword               = u32
type DataTypeDword32             = u64
type DataTypeDword64             = u64
type DataTypeDwordLong           = u64
type DataTypeFloat               = f32
type DataTypeHalfPtr             = i16
type DataTypeHFile               = int
type DataTypeHResult             = i64
type DataTypeInt                 = int
type DataTypeInt8                = i8
type DataTypeInt16               = i16
type DataTypeInt32               = int
type DataTypeInt64               = i64
type DataTypeIntPtr              = int
type DataTypeLong                = i64
type DataTypeLong32              = int
type DataTypeLong64              = i64
type DataTypeLongLong            = i64
type DataTypeLongPtr             = i64
type DataTypeLParam              = u64
type DataTypeLPByte              = u64
type DataTypeLPBool              = u64
type DataTypeLPColorRef          = u64
type DataTypeLPCStr              = u64
type DataTypeLPCTStr             = u64
type DataTypeLPCVoid             = u64
type DataTypeLPCWStr             = u64
type DataTypePInt                = int
type DataTypeLPInt               = u64
type DataTypeLPLong              = u64
type DataTypeLPTStr              = u64
type DataTypeLPVoid              = u64
type DataTypeLPWord              = u64
type DataTypeLPWStr              = u64
type DataTypePBool               = u32
type DataTypePBoolean            = u32
type DataTypePByte               = u32
type DataTypePChar               = u32
type DataTypePCStr               = u32
type DataTypePCTStr              = u32
type DataTypePCWStr              = u32
type DataTypePDword              = u32
type DataTypePDword32            = u32
type DataTypePDword64            = u32
type DataTypePDwordLong          = u32
type DataTypePDwordPtr           = u32
type DataTypePFloat              = u32
type DataTypePHalfPtr            = u32
type DataTypePHandle             = u32
type DataTypePHKey               = u32
type DataTypePInt8               = u32
type DataTypePInt16              = u32
type DataTypePInt32              = u32
type DataTypePInt64              = u32
type DataTypePIntPtr             = u32
type DataTypePLcID               = u32
type DataTypePLong               = u32
type DataTypePLong32             = u32
type DataTypePLong64             = u32
type DataTypePLongLong           = u32
type DataTypePLongPtr            = u32
type DataTypePointer32           = u32
type DataTypePointer64           = u64
type DataTypePointerSigned       = int
type DataTypePointerUnsigned     = u32
type DataTypePShort              = u32
type DataTypePSizeT              = u32
type DataTypePSSizeT             = u32
type DataTypePStr                = u32
type DataTypePTByte              = u32
type DataTypePTChar              = u32
type DataTypePTStr               = u32
type DataTypePWChar              = u32
type DataTypePWord               = u32
type DataTypePWStr               = u32
type DataTypePUChar              = u32
type DataTypePUHalfPtr           = u32
type DataTypePUInt               = u32
type DataTypePUInt8              = u32
type DataTypePUInt16             = u32
type DataTypePUInt32             = u32
type DataTypePUInt64             = u32
type DataTypePUIntPtr            = u32
type DataTypePULong              = u32
type DataTypePULong32            = u32
type DataTypePULong64            = u32
type DataTypePULongLong          = u32
type DataTypePULongPtr           = u32
type DataTypePUShort             = u32
type DataTypePVoid               = u32
type DataTypeQWord               = i64
type DataTypeShort               = i16
type DataTypeUChar               = u8
type DataTypeUHalfPtr            = u16
type DataTypeUInt                = u32
type DataTypeUInt8               = u8
type DataTypeUInt16              = u16
type DataTypeUInt32              = u32
type DataTypeUInt64              = u64
type DataTypeUIntPtr             = u32
type DataTypeULong               = u64
type DataTypeULong32             = u32
type DataTypeULong64             = u64
type DataTypeULongLong           = u64
type DataTypeULongPtr            = u64
type DataTypeUnicodeString       = string
type DataTypeUShort              = u16
// type DataTypeVoid                = any
type DataTypeWChar               = rune
type DataTypeWord                = u16

type DataTypeAtom                = u16   // DataTypeWord
type DataTypeBoolean             = u8    // DataTypeByte
type DataTypeChar                = i8    // DataTypeCChar
type DataTypeColorRef            = u32   // DataTypeDword
type DataTypeDwordPtr            = u64   // DataTypeUlongPtr
type DataTypeHandle              = u32   // DataTypePVoid
type DataTypeLangID              = u32   // DataTypeDword
type DataTypeLcID                = u32   // DataTypeDword
type DataTypeLcType              = u32   // DataTypeDword
type DataTypeLGrpID              = u32   // DataTypeDword
type DataTypeLResult             = u64   // DataTypeLongPtr
type DataTypeSCLock              = u32   // DataTypeLPVoid
type DataTypeSizeT               = u64   // DataTypeULongPtr
type DataTypeSSizeT              = i64   // DataTypeLongPtr
type DataTypeTByte               = rune  // DataTypeWChar
type DataTypeTChar               = rune  // DataTypeWChar
type DataTypeUSN                 = i64   // DataTypeLongLong
type DataTypeWParam              = u32   // DataTypeUIntPtr

type DataTypeHAccel              = u32   // DataTypeHandle
type DataTypeHBitmap             = u32   // DataTypeHandle
type DataTypeHBrush              = u32   // DataTypeHandle
type DataTypeHColorSpace         = u32   // DataTypeHandle
type DataTypeHConv               = u32   // DataTypeHandle
type DataTypeHConvList           = u32   // DataTypeHandle
type DataTypeHDC                 = u32   // DataTypeHandle
type DataTypeHDDEData            = u32   // DataTypeHandle
type DataTypeHDesk               = u32   // DataTypeHandle
type DataTypeHDrop               = u32   // DataTypeHandle
type DataTypeHDwp                = u32   // DataTypeHandle
type DataTypeHEnhMetafile        = u32   // DataTypeHandle
type DataTypeHFont               = u32   // DataTypeHandle
type DataTypeHGDIObj             = u32   // DataTypeHandle
type DataTypeHGlobal             = u32   // DataTypeHandle
type DataTypeHHook               = u32   // DataTypeHandle
type DataTypeHIcon               = u32   // DataTypeHandle
type DataTypeHInstance           = u32   // DataTypeHandle
type DataTypeHKey                = u32   // DataTypeHandle
type DataTypeHKL                 = u32   // DataTypeHandle
type DataTypeHLocal              = u32   // DataTypeHandle
type DataTypeHLPHandle           = u32   // DataTypeHandle
type DataTypeHMenu               = u32   // DataTypeHandle
type DataTypeHMetafile           = u32   // DataTypeHandle
type DataTypeHMonitor            = u32   // DataTypeHandle
type DataTypeHPalette            = u32   // DataTypeHandle
type DataTypeHPen                = u32   // DataTypeHandle
type DataTypeHRg                 = u32   // DataTypeHandle
type DataTypeHRsrc               = u32   // DataTypeHandle
type DataTypeHSZ                 = u32   // DataTypeHandle
type DataTypeHWinsta             = u32   // DataTypeHandle
type DataTypeHWnd                = u32   // DataTypeHandle
type DataTypeSCHandle            = u32   // DataTypeHandle
type DataTypeServiceStatusHandle = u32   // DataTypeHandle

type DataTypeHCursor             = u32   // DataTypeHIcon
type DataTypeHModule             = u32   // DataTypeHInstance
