module main

fn main() {
	println("${project_name} ${version}")
}
