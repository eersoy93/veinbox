/* DESCRIPTION: VeinBox simulation constants source file
 * AUTHOR: Erdem Ersoy (eersoy93)
 * See README.md for copyright and license.
 */

module simulation

const is_unicode = true
const is_win_64  = false
const win_ver    = u32(0x0502)
