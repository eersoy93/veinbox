/* DESCRIPTION: VeinBox simulation data types source file
 * AUTHOR: Erdem Ersoy (eersoy93)
 * See README.md for copyright and license.
 */

module simulation

type DataTypeBool            = int
type DataTypeByte            = u8
type DataTypeCChar           = i8
type DataTypeDword           = u32
type DataTypeDword32         = u64
type DataTypeDword64         = u64
type DataTypeDwordLong       = u64
type DataTypeFloat           = f32
type DataTypeHalfPtr         = i16
type DataTypeHFile           = int
type DataTypeHResult         = i64
type DataTypeInt             = int
type DataTypeInt8            = i8
type DataTypeInt16           = i16
type DataTypeInt32           = int
type DataTypeInt64           = i64
type DataTypeIntPtr          = int
type DataTypeLong            = i64
type DataTypeLong32          = int
type DataTypeLong64          = i64
type DataTypeLongLong        = i64
type DataTypeLongPtr         = i64
type DataTypeLPBool          = bool
type DataTypeLPInt           = int
type DataTypeLPLong          = i64
type DataTypeLPVoid          = u32
type DataTypeLPCStr          = u32
type DataTypeLPCVoid         = u32
type DataTypePInt            = int
type DataTypePointer32       = u32
type DataTypePointer64       = u64
type DataTypePointerSigned   = u32
type DataTypePointerUnsigned = u32
type DataTypePVoid           = u32
type DataTypeQWord           = i64
type DataTypeShort           = i16
type DataTypeUChar           = u8
type DataTypeUHalfPtr        = u16
type DataTypeUInt            = u32
type DataTypeUInt8           = u8
type DataTypeUInt16          = u16
type DataTypeUInt32          = u32
type DataTypeUInt64          = u64
type DataTypeUIntPtr         = u32
type DataTypeULong           = u64
type DataTypeULong32         = u32
type DataTypeULong64         = u64
type DataTypeULongLong       = u64
type DataTypeULongPtr        = u64
type DataTypeUnicodeString   = string
type DataTypeUShort          = u16
type DataTypeWChar           = rune
type DataTypeWord            = u16
// type DataTypeVoid          = any

type DataTypeAtom       = u16   // DataTypeWord
type DataTypeBoolean    = u8    // DataTypeByte
type DataTypeChar       = i8    // DataTypeCChar
type DataTypeColorRef   = u32   // DataTypeDword
type DataTypeDwordPtr   = u64   // DataTypeUlongPtr
type DataTypeHandle     = u32   // DataTypePVoid
type DataTypeLangID     = u32   // DataTypeDword
type DataTypeLcID       = u32   // DataTypeDword
type DataTypeLcType     = u32   // DataTypeDword
type DataTypeLGrpID     = u32   // DataTypeDword
type DataTypeLParam     = i64   // DataTypeLongPtr
type DataTypeLPByte     = u8    // DataTypeByte
type DataTypeLPColorRef = u32   // DataTypeDword
type DataTypeLPCWStr    = rune  // DataTypeWChar
type DataTypeLPWord     = u16   // DataTypeWord
type DataTypeLPWStr     = rune  // DataTypewChar
type DataTypeLResult    = u64   // DataTypeLongPtr
type DataTypePBool      = int   // DataTypeBool
type DataTypePByte      = u8    // DataTypeByte
type DataTypePChar      = i8    // DataTypeChar
type DataTypePCStr      = i8    // DataTypeChar
type DataTypePCWStr     = rune  // DataTypeWChar
type DataTypePDword     = u32   // DataTypeDword
type DataTypePDwordLong = u64   // DataTypeDwordLong
type DataTypePFloat     = f32   // DataTypeFloat
type DataTypePHalfPtr   = i16   // DataTypeHalfPtr
type DataTypePInt8      = i8    // DataTypeInt8
type DataTypePInt16     = i16   // DataTypeInt16
type DataTypePInt32     = int   // DataTypeInt32
type DataTypePInt64     = i64   // DataTypeInt64
type DataTypePIntPtr    = int   // DataTypeIntPtr
type DataTypePLong      = i64   // DataTypeLong
type DataTypePLong32    = int   // DataTypeLong32
type DataTypePLong64    = i64   // DataTypeLong64
type DataTypePLongLong  = i64   // DataTypeLongLong
type DataTypePLongPtr   = i64   // DataTypeLongPtr
type DataTypePShort     = i16   // DataTypeShort
type DataTypePUChar     = u8    // DataTypeUChar
type DataTypePUHalfPtr  = u16   // DataTypeUHalfPtr
type DataTypePUInt      = u32   // DataTypeUInt
type DataTypePUInt8     = u8    // DataTypeUInt8
type DataTypePUInt16    = u16   // DataTypeUInt16
type DataTypePUInt32    = u32   // DataTypeUInt32
type DataTypePUInt64    = u64   // DataTypeUInt64
type DataTypePUIntPtr   = u32   // DataTypeUIntPtr
type DataTypePULong     = u64   // DataTypeULong
type DataTypePULong32   = u32   // DataTypeULong32
type DataTypePULong64   = u64   // DataTypeULong64
type DataTypePULongLong = u64   // DataTypeULongLong
type DataTypePULongPtr  = u64   // DataTypeULongPtr
type DataTypePUShort    = u16   // DataTypeUShort
type DataTypePWChar     = rune  // DataTypeWChar
type DataTypePWord      = u16   // DataTypeWord
type DataTypePWStr      = rune  // DataTypeWChar
type DataTypeSCLock     = u32   // DataTypeLPVoid
type DataTypeSizeT      = u64   // DataTypeULongPtr
type DataTypeSSizeT     = i64   // DataTypeLongPtr
type DataTypeTByte      = rune  // DataTypeWChar
type DataTypeTChar      = rune  // DataTypeWChar
type DataTypeUSN        = i64   // DataTypeLongLong
type DataTypeWParam     = u32   // DataTypeUIntPtr

type DataTypeHAccel              = u32   // DataTypeHandle
type DataTypeHBitmap             = u32   // DataTypeHandle
type DataTypeHBrush              = u32   // DataTypeHandle
type DataTypeHColorSpace         = u32   // DataTypeHandle
type DataTypeHConv               = u32   // DataTypeHandle
type DataTypeHConvList           = u32   // DataTypeHandle
type DataTypeHDC                 = u32   // DataTypeHandle
type DataTypeHDDEData            = u32   // DataTypeHandle
type DataTypeHDesk               = u32   // DataTypeHandle
type DataTypeHDrop               = u32   // DataTypeHandle
type DataTypeHDwp                = u32   // DataTypeHandle
type DataTypeHEnhMetafile        = u32   // DataTypeHandle
type DataTypeHFont               = u32   // DataTypeHandle
type DataTypeHGDIObj             = u32   // DataTypeHandle
type DataTypeHGlobal             = u32   // DataTypeHandle
type DataTypeHHook               = u32   // DataTypeHandle
type DataTypeHIcon               = u32   // DataTypeHandle
type DataTypeHInstance           = u32   // DataTypeHandle
type DataTypeHKey                = u32   // DataTypeHandle
type DataTypeHKL                 = u32   // DataTypeHandle
type DataTypeHLocal              = u32   // DataTypeHandle
type DataTypeHLPHandle           = u32   // DataTypeHandle
type DataTypeHMenu               = u32   // DataTypeHandle
type DataTypeHMetafile           = u32   // DataTypeHandle
type DataTypeHMonitor            = u32   // DataTypeHandle
type DataTypeHPalette            = u32   // DataTypeHandle
type DataTypeHPen                = u32   // DataTypeHandle
type DataTypeHRg                 = u32   // DataTypeHandle
type DataTypeHRsrc               = u32   // DataTypeHandle
type DataTypeHSZ                 = u32   // DataTypeHandle
type DataTypeHWinsta             = u32   // DataTypeHandle
type DataTypeHWnd                = u32   // DataTypeHandle
type DataTypeLPCTStr             = rune  // DataTypeLPCWStr
type DataTypeLPTStr              = rune  // DataTypeLPWStr
type DataTypePBoolean            = u8    // DataTypeBoolean
type DataTypePCTStr              = u32   // DataTypeWChar
type DataTypePDword32            = u64   // DataTypePDword
type DataTypePDword64            = u64   // DataTypePDword
type DataTypePDwordPtr           = u64   // DataTypeDwordPtr
type DataTypePHandle             = u32   // DataTypeHandle
type DataTypePLcID               = u32   // DataTypeLcID
type DataTypePSizeT              = u64   // DataTypeSizeT
type DataTypePSSizeT             = i64   // DataTypeSSizeT
type DataTypePStr                = i8    // DataTypeChar
type DataTypePTByte              = rune  // DataTypeTByte
type DataTypePTChar              = rune  // DataTypeTChar
type DataTypePTStr               = rune  // DataTypeLPWStr
type DataTypeSCHandle            = u32   // DataTypeHandle
type DataTypeServiceStatusHandle = u32   // DataTypeHandle

type DataTypeHCursor      = u32   // DataTypeHIcon
type DataTypeHModule      = u32   // DataTypeHInstance
type DataTypePHKey        = u32   // DataTypeHKey
