/* DESCRIPTION: VeinBox main source file
 * AUTHOR: Erdem Ersoy (eersoy93)
 * See README.md for copyright and license.
 */

module main

fn main() {
	println("${project_name} ${version}")
}
