module main

const project_name   = "VeinBox"

const version_major  = u8(0)
const version_middle = u8(0)
const version_minor  = u8(1)

const version        = "${version_major}.${version_middle}.${version_minor}"
