/* DESCRIPTION: VeinBox simulation data types source file
 * AUTHOR: Erdem Ersoy (eersoy93)
 * See README.md for copyright and license.
 */

module simulation

type DataTypeBool          = bool
type DataTypeByte          = u8
type DataTypeCChar         = i8
type DataTypeDword         = u32
type DataTypeDword32       = u64
type DataTypeDword64       = u64
type DataTypeDwordLong     = u64
type DataTypeFloat         = f32
type DataTypeHalfPtr       = i16
type DataTypeHFile         = int
type DataTypeHResult       = i64
type DataTypeInt           = int
type DataTypeInt8          = i8
type DataTypeInt16         = i16
type DataTypeInt32         = int
type DataTypeInt64         = i64
type DataTypeIntPtr        = int
type DataTypeLong          = i64
type DataTypeLong32        = int
type DataTypeLong64        = i64
type DataTypeLongLong      = i64
type DataTypeLongPtr       = i64
type DataTypeLPBool        = bool
type DataTypeLPInt         = int
type DataTypeLPLong        = i64
type DataTypeLPVoid        = u32
type DataTypeLPCStr        = u32
type DataTypeLPCVoid       = u32
type DataTypePVoid         = u32
type DataTypeUChar         = u8
type DataTypeUHalfPtr      = u16
type DataTypeUInt          = u32
type DataTypeUInt8         = u8
type DataTypeUInt16        = u16
type DataTypeUInt32        = u32
type DataTypeUInt64        = u64
type DataTypeUIntPtr       = u32
type DataTypeULong         = u64
type DataTypeULong32       = u32
type DataTypeULong64       = u64
type DataTypeULongLong     = u64
type DataTypeULongPtr      = u64
type DataTypeUnicodeString = string
type DataTypeUShort        = u16
type DataTypeWChar         = rune
type DataTypeWord          = u16
// type DataTypeVoid          = any

type DataTypeAtom       = DataTypeWord
type DataTypeBoolean    = DataTypeByte
type DataTypeChar       = DataTypeCChar
type DataTypeColorRef   = DataTypeDword
type DataTypeDwordPtr   = DataTypeUlongPtr
type DataTypeHandle     = DataTypePVoid
type DataTypeLangID     = DataTypeDword
type DataTypeLcID       = DataTypeDword
type DataTypeLcType     = DataTypeDword
type DataTypeLGrpID     = DataTypeDword
type DataTypeLParam     = DataTypeLongPtr
type DataTypeLPByte     = DataTypeByte
type DataTypeLPColorRef = DataTypeDword
type DataTypeLPCWStr    = DataTypeWChar
type DataTypeLPWord     = DataTypeWord
type DataTypeLPWStr     = DataTypewChar
type DataTypeLResult    = DataTypeLongPtr
type DataTypePBool      = DataTypeBool
type DataTypePBoolean   = DataTypeBoolean
type DataTypePByte      = DataTypeByte
type DataTypePChar      = DataTypeChar
type DataTypePCStr      = DataTypeChar
type DataTypePCWStr     = DataTypeWChar
type DataTypeTByte      = DataTypeWChar
type DataTypeTChar      = DataTypeWChar
type DataTypeUSN        = DataTypeLongLong
type DataTypeWParam     = DataTypeUIntPtr

type DataTypeHAccel       = DataTypeHandle
type DataTypeHBitmap      = DataTypeHandle
type DataTypeHBrush       = DataTypeHandle
type DataTypeHColorSpace  = DataTypeHandle
type DataTypeHConv        = DataTypeHandle
type DataTypeHConvList    = DataTypeHandle
type DataTypeHDC          = DataTypeHandle
type DataTypeHDDEData     = DataTypeHandle
type DataTypeHDesk        = DataTypeHandle
type DataTypeHDrop        = DataTypeHandle
type DataTypeHDwp         = DataTypeHandle
type DataTypeHEnhMetafile = DataTypeHandle
type DataTypeHFont        = DataTypeHandle
type DataTypeHGDIObj      = DataTypeHandle
type DataTypeHGlobal      = DataTypeHandle
type DataTypeHHook        = DataTypeHandle
type DataTypeHIcon        = DataTypeHandle
type DataTypeHInstance    = DataTypeHandle
type DataTypeHKey         = DataTypeHandle
type DataTypeHKL          = DataTypeHandle
type DataTypeHLocal       = DataTypeHandle
type DataTypeHLPHandle    = DataTypeHandle
type DataTypeHMenu        = DataTypeHandle
type DataTypeHMetafile    = DataTypeHandle
type DataTypeHMonitor     = DataTypeHandle
type DataTypeHPalette     = DataTypeHandle
type DataTypeHPen         = DataTypeHandle
type DataTypeHRg          = DataTypeHandle
type DataTypeHRsrc        = DataTypeHandle
type DataTypeHSZ          = DataTypeHandle
type DataTypeHWinsta      = DataTypeHandle
type DataTypeHWnd         = DataTypeHandle
type DataTypeLPCTStr      = DataTypeLPCWStr
type DataTypeLPTStr       = DataTypeLPWStr
type DataTypePCTStr       = DataTypeWChar

type DataTypeHCursor      = DataTypeHIcon
type DataTypeHModule      = DataTypeHInstance
